package yapp_pkg;

  // import the UVM library
  import uvm_pkg::*;

  // include the UVM macros
  `include "uvm_macros.svh"

  // include the YAPP packet definition
  `include "yapp_packet.sv" 
  `include  "yapp_tx_monitor.sv"
  `include  "yapp_tx_sequencer.sv"
  `include  "yapp_tx_seqs.sv"
  `include  "yapp_tx_driver.sv"
  `include  "yapp_tx_agent.sv"
  `include  "yapp_tx_env.sv"
endpackage : yapp_pkg
